module cmp_unit(


);

endmodule